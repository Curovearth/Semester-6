module fa_df_19BEE0167(input a,b,cin,output sum,cout);
assign sum=a^b^cin;
assign cout=(a^b)&cin|(a&b);
endmodule
