

module ha_df_19BEE0167(input a,b,
			output sum,cout);
assign sum = a^b; 
assign cout = a&b; 
endmodule